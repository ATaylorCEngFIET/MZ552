library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package p_wave_Package is
    type t_sine_array is array (0 to 99) of std_logic_vector(15 downto 0);
    -- put python results below
    constant analog_wave : t_sine_array := (
        "0111111111111111",
        "1000100000001000",
        "1001000000001010",
        "1001011111111011",
        "1001111111010100",
        "1010011110001101",
        "1010111100011110",
        "1011011001111111",
        "1011110110101001",
        "1100010010010101",
        "1100101100111011",
        "1101000110010110",
        "1101011110011110",
        "1101110101001101",
        "1110001010011111",
        "1110011110001100",
        "1110110000010010",
        "1111000000101001",
        "1111001111010000",
        "1111011100000001",
        "1111100110111011",
        "1111101111111001",
        "1111110110111010",
        "1111111011111100",
        "1111111110111110",
        "1111111111111111",
        "1111111110111110",
        "1111111011111100",
        "1111110110111010",
        "1111101111111001",
        "1111100110111011",
        "1111011100000001",
        "1111001111010000",
        "1111000000101001",
        "1110110000010010",
        "1110011110001100",
        "1110001010011111",
        "1101110101001101",
        "1101011110011110",
        "1101000110010110",
        "1100101100111011",
        "1100010010010101",
        "1011110110101001",
        "1011011001111111",
        "1010111100011110",
        "1010011110001101",
        "1001111111010100",
        "1001011111111011",
        "1001000000001010",
        "1000100000001000",
        "0111111111111111",
        "0111011111110110",
        "0110111111110100",
        "0110100000000011",
        "0110000000101010",
        "0101100001110001",
        "0101000011100000",
        "0100100101111111",
        "0100001001010101",
        "0011101101101001",
        "0011010011000011",
        "0010111001101000",
        "0010100001100000",
        "0010001010110001",
        "0001110101011111",
        "0001100001110010",
        "0001001111101100",
        "0000111111010101",
        "0000110000101110",
        "0000100011111101",
        "0000011001000011",
        "0000010000000101",
        "0000001001000100",
        "0000000100000010",
        "0000000001000000",
        "0000000000000000",
        "0000000001000000",
        "0000000100000010",
        "0000001001000100",
        "0000010000000101",
        "0000011001000011",
        "0000100011111101",
        "0000110000101110",
        "0000111111010101",
        "0001001111101100",
        "0001100001110010",
        "0001110101011111",
        "0010001010110001",
        "0010100001100000",
        "0010111001101000",
        "0011010011000011",
        "0011101101101001",
        "0100001001010101",
        "0100100101111111",
        "0101000011100000",
        "0101100001110001",
        "0110000000101010",
        "0110100000000011",
        "0110111111110100",
        "0111011111110110"
    );
end p_wave_Package;